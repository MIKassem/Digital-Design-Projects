
module ALU_tb;
  reg [3:0] C;
  reg [7:0] A, B;
  wire [7:0] s;
  wire cout;
  ALU uut (C,A,B,s,cout);

initial begin
  $dumpfile("waf.vcd");
  $dumpvars(1);
A = 8'b00000000;B = 8'b11111110; C=4'b0001;
#10 A = 8'b00110010;B = 8'b00110010; C = 4'b0001;
#10 A = 8'b00110010;B = 8'b01001011; C = 4'b0001;
#10 A = 8'b11001110;B = 8'b10110101; C = 4'b0001;
#10 A = 8'b01100100;B = 8'b10011100; C = 4'b0001;
  
  
#10 A = 8'b00000000;B = 8'b11111110; C=4'b0010;
#10 A = 8'b00110010;B = 8'b00110010; C = 4'b0010;
#10 A = 8'b00110010;B = 8'b01001011; C = 4'b0010;
#10 A = 8'b11001110;B = 8'b10110101; C = 4'b0010;
#10 A = 8'b01100100;B = 8'b10011100; C = 4'b0010;
  
  
#10 A = 8'b00000000;B = 8'b11111110; C=4'b0011;
#10 A = 8'b00110010;B = 8'b00110010; C = 4'b0011;
#10 A = 8'b00110010;B = 8'b01001011; C = 4'b0011;
#10 A = 8'b11001110;B = 8'b10110101; C = 4'b0011;
#10 A = 8'b01100100;B = 8'b10011100; C = 4'b0011;


#10 A = 8'b00000000;B = 8'b11111110; C=4'b0100;
#10 A = 8'b00110010;B = 8'b00110010; C = 4'b0100;
#10 A = 8'b00110010;B = 8'b01001011; C = 4'b0100;
#10 A = 8'b11001110;B = 8'b10110101; C = 4'b0100;
#10 A = 8'b01100100;B = 8'b10011100; C = 4'b0100;

  
#10 A = 8'b00000000;B = 8'b11111110; C=4'b0110;
#10 A = 8'b00110010;B = 8'b00110010; C = 4'b0110;
#10 A = 8'b00110010;B = 8'b01001011; C = 4'b0110;
#10 A = 8'b11001110;B = 8'b10110101; C = 4'b0110;
#10 A = 8'b01100100;B = 8'b10011100; C = 4'b0110;

  
#10 A = 8'b00000000;B = 8'b11111110; C=4'b0111;
#10 A = 8'b00110010;B = 8'b00110010; C = 4'b0111;
#10 A = 8'b00110010;B = 8'b01001011; C = 4'b0111;
#10 A = 8'b11001110;B = 8'b10110101; C = 4'b0111;
#10 A = 8'b01100100;B = 8'b10011100; C = 4'b0111;
  
#10 A = 8'b11001101; C = 4'b1000;
#10 A = 8'b01010101; C = 4'b1000;
#10 A = 8'b11001101; C = 4'b1000;
#10 A = 8'b01010101; C = 4'b1000;

#10 A = 8'b11001101; C = 4'b1001;
#10 A = 8'b01010101; C = 4'b1001;
#10 A = 8'b11001101; C = 4'b1001;
#10 A = 8'b01010101; C = 4'b1001;
  
#10 A = 8'b11001101; C = 4'b1010;
#10 A = 8'b01010101; C = 4'b1010;
#10 A = 8'b11001101; C = 4'b1010;
#10 A = 8'b01010101; C = 4'b1010;
  
#10 A = 8'b11001101; C = 4'b1011;
#10 A = 8'b01010101; C = 4'b1011;
#10 A = 8'b11001101; C = 4'b1011;
#10 A = 8'b01010101; C = 4'b1011;
  
#10 A = 8'b11001101; C = 4'b1100;
#10 A = 8'b01010101; C = 4'b1100;
#10 A = 8'b11001101; C = 4'b1100;
#10 A = 8'b01010101; C = 4'b1100;

  
#10 A = 8'b11001101; C = 4'b1101;
#10 A = 8'b01010101; C = 4'b1101;
#10 A = 8'b11001101; C = 4'b1101;
#10 A = 8'b01010101; C = 4'b1101;
  
end
endmodule